module types

pub struct Image {
pub:
	id string [json: Id]
}
